module FLAGS
(
    
);
endmodule