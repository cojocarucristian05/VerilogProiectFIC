module CPU
(

);

endmodule