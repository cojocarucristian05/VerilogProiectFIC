module STACK
(

);
endmodule