module REGISTERS
(

);
endmodule