module FLAGS
(

);
endmodule